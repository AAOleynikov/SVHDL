-------------------------------------------------------------------------------
--
-- Title       : 
-- Design      : lab4
-- Author      : 666anton2005xr@gmail.com
-- Company     : 666anton2005xr@gmail.com
--
-------------------------------------------------------------------------------
--
-- File        : jk_with_polar_control_TB.vhd
-- Generated   : Sun May  5 19:22:55 2024
-- From        : C:\Users\666an\Documents\BMSTU\MVHDL\Labs (2)\lab4\src\WAVES\jk_with_polar_control_TB_settings.txt
-- By          : tb_generator.pl ver. ver 1.2s
--
-------------------------------------------------------------------------------
--
-- Description : declaration of TEST_PINS package
--
-------------------------------------------------------------------------------
--The TEST_PINS package contains declaration of enumerated type named TEST_PINS.
--This declaration contains one enumerated value for each port
-- find in test vector file:
--An order of declared values match the order of ports in test vector file.

package UUT_TEST_PINS is
type TEST_PINS is (
--The test vector file:  does not contains any test vectors for the port of the UUT: jk_with_polar_control,
--therefore the TEST_PINS type has no elements and causes compilation error.
);
end UUT_TEST_PINS;
